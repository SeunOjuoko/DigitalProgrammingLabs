module Lab4(clk,temp,select,disp_drive,temp0,temp1,temp2,temp3,avg);
	// includes the display drivers
	input clk;
	input [9:0] temp;
	input [3:0] select;
	output [20:0] disp_drive;
	
	output [9:0] avg,temp0,temp1,temp2,temp3;
	
	reg [9:0] temp0,temp1,temp2,temp3;//outputs to decoder
	reg [11:0] sum1;
	reg [9:0] avg;
	wire[9:0] avg1;
	assign avg1=avg;

	bcd_decode_display b1(clk,avg,disp_drive);
	always @(posedge clk)
		begin
			case (select)
				4'b1110 : temp0 = temp; // segments lit
				4'b1101 : temp1 = temp;
				4'b1011 : temp2 = temp;
				4'b0111 : temp3 = temp;
				default :;
				endcase
			sum1=temp0+temp1+temp2+temp3;
			avg=sum1/4;
	end
endmodule

module bcd_decode_display(clk,number,disp_drive);
	// includes the display drivers
	input clk;
	input [9:0] number;
	output [20:0] disp_drive;//outputs to display segments
	reg [3:0] numb_bcd0,numb_bcd1,numb_bcd2;
	wire [3:0] n1,n2,n3;
	assign n1 = numb_bcd0;
	assign n2 = numb_bcd1;
	assign n3 = numb_bcd2;
	// instantiate each display driver
	display_drv units(clk,n1,disp_drive[6:0]); // Least significant digit
	display_drv tenths(clk,n2,disp_drive[13:7]);
	display_drv hundredths(clk,n2,disp_drive[20:14]);
	// bcd conversion units, tens and hundreds
	always @(posedge clk)
		begin
		numb_bcd2 = number/100;
		numb_bcd1 = (number%100)/10;
		numb_bcd0 = (number%100)%10;
	end
endmodule

module display_drv(clk,number,display);
	input clk;
	input [3:0] number;
	output [6:0] display;
	reg [6:0] d;
	assign display = d; // active high
	// on clock edge update display
	always @(posedge clk )
		begin
		if (number < 10)
			begin
				case (number)
				4'd0 : d <= 7'b1000000; // segments lit
				4'd1 : d <= 7'b1111001;
				4'd2 : d <= 7'b0100100;
				4'd3 : d <= 7'b0110000;
				4'd4 : d <= 7'b0011001;
				4'd5 : d <= 7'b0010010;
				4'd6 : d <= 7'b0000010;
				4'd7 : d <= 7'b1111000;
				4'd8 : d <= 7'b0000000;
				4'd9 : d <= 7'b0011000;
				default : d <= 7'b1111111; // off
				endcase
			end
		else d <= 7'b0001110; // 'F'	
	end
endmodule
